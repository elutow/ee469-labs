// Writes back the result of executor to the regfile

module regfilewriter(
        input wire clk,
        input wire nreset,
        input logic enable,
        output logic ready
    );
endmodule
