`ifndef _CPU_CONSTANTS_SVH_
`define _CPU_CONSTANTS_SVH_

// TODO: Move macros to include
// Register & instruction depths
`define BIT_WIDTH 32
// Size of register file
`define REG_COUNT 16
// TODO: Change to correct number of instructions
`define INST_COUNT 64
// DEBUG_BYTES Must be power of 2
`define DEBUG_BYTES 32

`endif
